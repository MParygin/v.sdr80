`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: makkosik
// 
// Create Date:    14:51:10 02/16/2012 
// Design Name: 
// Module Name:    sincos 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description:    Sin Cos Lut (17 bits)
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sincos(
    input wire clk,
	 input wire [11:0] phase,
	 output reg [16:0] out_sin,
	 output reg [16:0] out_cos
);

// quadrant
wire [1:0] quadrant_sin = phase[11:10];
wire [1:0] quadrant_cos = phase[11:10];

// virtual address sin
wire [9:0] vaddr_sin = (quadrant_sin[0] == 1'b0) ? phase[9:0] : ~phase[9:0];
wire [9:0] vaddr_cos = (quadrant_cos[0] == 1'b0) ? phase[9:0] : ~phase[9:0];


// LUT
wire [15:0] sin_out;
wire [15:0] cos_out;
RAMB16_S18_S18 #(
.INIT_00(256'h061605B1054D04E80484041F03BB035602F1028D022801C4015F00FB00960032),
.INIT_01(256'h0C5D0BF90B940B300ACB0A670A02099E093908D50871080C07A8074306DF067A),
.INIT_02(256'h12A2123E11DA1176111110AD10490FE40F800F1C0EB70E530DEF0D8A0D260CC1),
.INIT_03(256'h18E51881181D17B9175516F1168D162815C4156014FC1498143313CF136B1307),
.INIT_04(256'h1F241EC01E5C1DF81D951D311CCD1C691C051BA11B3D1AD91A751A1119AD1949),
.INIT_05(256'h255E24FA2497243323D0236C230922A5224221DE217A211720B3204F1FEB1F88),
.INIT_06(256'h2B922B2F2ACC2A692A0629A2293F28DC2879281627B2274F26EC2688262525C1),
.INIT_07(256'h31C0315D30FA309830352FD22F6F2F0D2EAA2E472DE42D812D1E2CBB2C582BF5),
.INIT_08(256'h37E53783372136BF365D35FB3598353634D43471340F33AC334A32E732853222),
.INIT_09(256'h3E033DA13D403CDE3C7C3C1B3BB93B573AF53A933A3139D0396E390C38AA3848),
.INIT_0A(256'h441643B5435442F34292423141D0416F410E40AD404B3FEA3F893F273EC63E64),
.INIT_0B(256'h4A1F49BF495F48FF489E483E47DD477D471C46BC465B45FA459A453944D84477),
.INIT_0C(256'h501D4FBE4F5E4EFF4E9F4E3F4DDF4D804D204CC04C604C004BA04B404AE04A80),
.INIT_0D(256'h560F55B0555154F25493543553D65377531752B8525951FA519B513B50DC507D),
.INIT_0E(256'h5BF35B955B375AD95A7B5A1D59BF5961590258A4584657E75789572A56CC566D),
.INIT_0F(256'h61C9616C610F60B260545FF75F9A5F3D5EDF5E825E255DC75D6A5D0C5CAE5C50),
.INIT_10(256'h678F673366D7667B661F65C36567650A64AE645163F56398633C62DF62826225),
.INIT_11(256'h6D466CEB6C906C356BDA6B7F6B246AC86A6D6A1169B6695A68FF68A3684767EB),
.INIT_12(256'h72EC7292723971DF7184712A70D07076701B6FC16F676F0C6EB16E576DFC6DA1),
.INIT_13(256'h7881782877CF7776771D76C4766B761275B9755F750674AD745373FA73A07346),
.INIT_14(256'h7E027DAB7D537CFB7CA47C4C7BF47B9C7B447AEC7A937A3B79E3798A793278D9),
.INIT_15(256'h8371831A82C4826D821781C0816A811380BC8065800E7FB77F607F097EB17E5A),
.INIT_16(256'h88CB8876882187CB8776872186CB8676862085CB8575851F84C98473841D83C7),
.INIT_17(256'h8E108DBC8D688D148CC08C6C8C188BC48B708B1B8AC78A728A1E89C989748920),
.INIT_18(256'h933F92EC929A924791F591A2915090FD90AA905790048FB18F5D8F0A8EB78E63),
.INIT_19(256'h9857980697B59764971396C29670961F95CE957C952A94D99487943593E39391),
.INIT_1A(256'h9D589D089CB99C699C1A9BCA9B7A9B2A9ADA9A8A9A3A99EA9999994998F898A8),
.INIT_1B(256'hA240A1F2A1A5A157A108A0BAA06CA01E9FCF9F809F329EE39E949E459DF69DA7),
.INIT_1C(256'hA710A6C4A677A62BA5DEA592A545A4F8A4ABA45EA411A3C4A376A329A2DCA28E),
.INIT_1D(256'hABC6AB7BAB30AAE5AA9BAA50AA04A9B9A96EA922A8D7A88BA840A7F4A7A8A75C),
.INIT_1E(256'hB061B018AFCFAF86AF3DAEF3AEAAAE60AE17ADCDAD83AD39ACEFACA5AC5AAC10),
.INIT_1F(256'hB4E1B49AB452B40BB3C3B37CB334B2ECB2A4B25CB214B1CCB183B13BB0F2B0AA),
.INIT_20(256'hB945B900B8BAB874B82FB7E9B7A3B75DB717B6D0B68AB643B5FDB5B6B56FB528),
.INIT_21(256'hBD8DBD49BD05BCC1BC7EBC39BBF5BBB1BB6DBB28BAE3BA9FBA5ABA15B9D0B98A),
.INIT_22(256'hC1B7C175C133C0F1C0AFC06DC02BBFE8BFA6BF63BF20BEDDBE9ABE57BE14BDD0),
.INIT_23(256'hC5C4C584C544C504C4C3C483C442C402C3C1C380C33FC2FEC2BDC27CC23AC1F9),
.INIT_24(256'hC9B2C974C936C8F7C8B9C87BC83CC7FDC7BEC780C740C701C6C2C683C643C603),
.INIT_25(256'hCD81CD45CD08CCCCCC90CC53CC17CBDACB9DCB60CB23CAE6CAA8CA6BCA2DC9EF),
.INIT_26(256'hD130D0F6D0BCD081D047D00CCFD2CF97CF5CCF21CEE6CEABCE6FCE34CDF8CDBC),
.INIT_27(256'hD4BFD487D44FD416D3DED3A6D36DD334D2FBD2C2D289D250D217D1DDD1A3D16A),
.INIT_28(256'hD82DD7F7D7C1D78BD754D71ED6E7D6B1D67AD643D60CD5D5D59DD566D52ED4F7),
.INIT_29(256'hDB7ADB46DB12DADEDAAADA75DA41DA0CD9D8D9A3D96ED939D903D8CED898D863),
.INIT_2A(256'hDEA5DE73DE41DE0FDDDDDDABDD79DD46DD13DCE1DCAEDC7BDC48DC14DBE1DBAD),
.INIT_2B(256'hE1ADE17EE14EE11EE0EEE0BEE08EE05EE02DDFFDDFCCDF9BDF6ADF39DF08DED6),
.INIT_2C(256'hE493E466E438E40BE3DDE3AFE381E353E325E2F6E2C8E299E26AE23BE20CE1DD),
.INIT_2D(256'hE756E72BE6FFE6D4E6A9E67DE651E625E5F9E5CDE5A0E574E547E51AE4EDE4C0),
.INIT_2E(256'hE9F5E9CCE9A3E97AE950E927E8FDE8D4E8AAE880E856E82BE801E7D6E7ACE781),
.INIT_2F(256'hEC70EC49EC22EBFBEBD4EBADEB86EB5EEB37EB0FEAE7EABFEA97EA6FEA46EA1E),
.INIT_30(256'hEEC6EEA2EE7DEE59EE34EE0FEDEAEDC5ED9FED7AED54ED2FED09ECE3ECBCEC96),
.INIT_31(256'hF0F8F0D6F0B3F091F06FF04CF029F006EFE3EFC0EF9DEF79EF56EF32EF0EEEEA),
.INIT_32(256'hF304F2E4F2C4F2A5F284F264F244F223F202F1E2F1C1F19FF17EF15DF13BF119),
.INIT_33(256'hF4EBF4CEF4B0F492F475F457F439F41BF3FCF3DEF3BFF3A0F381F362F343F324),
.INIT_34(256'hF6ACF691F676F65BF63FF624F608F5ECF5D0F5B4F598F57BF55FF542F525F508),
.INIT_35(256'hF847F82FF816F7FDF7E4F7CBF7B2F798F77EF765F74BF731F716F6FCF6E2F6C7),
.INIT_36(256'hF9BCF9A6F990F979F962F94CF935F91EF906F8EFF8D8F8C0F8A8F890F878F860),
.INIT_37(256'hFB0AFAF7FAE3FACFFABAFAA6FA92FA7DFA68FA53FA3EFA29FA13F9FEF9E8F9D2),
.INIT_38(256'hFC32FC21FC0FFBFEFBECFBDAFBC8FBB5FBA3FB91FB7EFB6BFB58FB45FB31FB1E),
.INIT_39(256'hFD33FD24FD15FD06FCF6FCE7FCD7FCC7FCB7FCA7FC97FC86FC76FC65FC54FC43),
.INIT_3A(256'hFE0CFE00FDF3FDE7FDDAFDCDFDBFFDB2FDA5FD97FD89FD7BFD6DFD5FFD50FD42),
.INIT_3B(256'hFEBFFEB5FEABFEA0FE96FE8BFE81FE76FE6BFE5FFE54FE48FE3DFE31FE25FE19),
.INIT_3C(256'hFF4AFF43FF3BFF33FF2BFF23FF1BFF12FF0AFF01FEF8FEEFFEE5FEDCFED3FEC9),
.INIT_3D(256'hFFAEFFA9FFA4FF9EFF99FF93FF8DFF87FF81FF7BFF74FF6EFF67FF60FF59FF52),
.INIT_3E(256'hFFEBFFE8FFE5FFE2FFDFFFDCFFD8FFD5FFD1FFCDFFC9FFC5FFC1FFBCFFB8FFB3),
.INIT_3F(256'hFFFFFFFFFFFFFFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF7FFF5FFF3FFF1FFEFFFED)
) RAM_Inst (
  .CLKA(clk),
  .CLKB(clk),
  .ENA(1'b1),
  .ENB(1'b1),
  .WEA(1'b0),
  .WEB(1'b0),
  .ADDRA(vaddr_sin),
  .ADDRB(vaddr_cos),
  .SSRA(1'b0),
  .SSRB(1'b0),
  .DIPA(2'b0),
  .DIPB(2'b0),
  .DOPA(),
  .DOPB(),
  .DIA(16'b0),
  .DIB(16'b0),
  .DOA(sin_out),
  .DOB(cos_out)
);

// temporary calcs
wire [16:0] tout_sin = {quadrant_sin[1], (quadrant_sin[1] == 1'b0) ? sin_out : ~sin_out + 1};
wire [16:0] tout_cos = {quadrant_sin[1], (quadrant_sin[1] == 1'b0) ? sin_out : ~sin_out + 1};

// reg assign
always @ (posedge clk)
begin
  out_sin <= tout_sin;
  out_cos <= tout_cos;
end

endmodule
